ilireset_inst : ilireset PORT MAP (
		data	 => data_sig,
		result	 => result_sig
	);
