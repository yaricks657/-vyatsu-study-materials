// megafunction wizard: %LPM_CLSHIFT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_clshift 

// ============================================================
// File Name: Shift1.v
// Megafunction Name(s):
// 			lpm_clshift
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.1 Build 350 03/24/2010 SP 2 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2010 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module Shift1 (
	data,
	distance,
	result);

	input	[16:0]  data;
	input	[1:0]  distance;
	output	[16:0]  result;

	wire [16:0] sub_wire0;
	wire  sub_wire1 = 1'h1;
	wire [16:0] result = sub_wire0[16:0];

	lpm_clshift	lpm_clshift_component (
				.distance (distance),
				.direction (sub_wire1),
				.data (data),
				.result (sub_wire0)
				// synopsys translate_off
				,
				.aclr (),
				.clken (),
				.clock (),
				.overflow (),
				.underflow ()
				// synopsys translate_on
				);
	defparam
		lpm_clshift_component.lpm_shifttype = "LOGICAL",
		lpm_clshift_component.lpm_type = "LPM_CLSHIFT",
		lpm_clshift_component.lpm_width = 17,
		lpm_clshift_component.lpm_widthdist = 2;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: PRIVATE: LPM_SHIFTTYPE NUMERIC "0"
// Retrieval info: PRIVATE: LPM_WIDTH NUMERIC "17"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: lpm_width_varies NUMERIC "0"
// Retrieval info: PRIVATE: lpm_widthdist NUMERIC "2"
// Retrieval info: PRIVATE: lpm_widthdist_style NUMERIC "1"
// Retrieval info: PRIVATE: port_direction NUMERIC "1"
// Retrieval info: CONSTANT: LPM_SHIFTTYPE STRING "LOGICAL"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_CLSHIFT"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "17"
// Retrieval info: CONSTANT: LPM_WIDTHDIST NUMERIC "2"
// Retrieval info: USED_PORT: data 0 0 17 0 INPUT NODEFVAL data[16..0]
// Retrieval info: USED_PORT: distance 0 0 2 0 INPUT NODEFVAL distance[1..0]
// Retrieval info: USED_PORT: result 0 0 17 0 OUTPUT NODEFVAL result[16..0]
// Retrieval info: CONNECT: @distance 0 0 2 0 distance 0 0 2 0
// Retrieval info: CONNECT: @data 0 0 17 0 data 0 0 17 0
// Retrieval info: CONNECT: result 0 0 17 0 @result 0 0 17 0
// Retrieval info: CONNECT: @direction 0 0 0 0 VCC 0 0 0 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift1.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift1.inc TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift1.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift1.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift1_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift1_bb.v TRUE
