-- megafunction wizard: %LPM_XOR%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: lpm_xor 

-- ============================================================
-- File Name: xor48.vhd
-- Megafunction Name(s):
-- 			lpm_xor
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 350 03/24/2010 SP 2 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY xor48 IS
	PORT
	(
		data		: IN STD_LOGIC_2D (47 DOWNTO 0, 47 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (47 DOWNTO 0)
	);
END xor48;


ARCHITECTURE SYN OF xor48 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (47 DOWNTO 0);

BEGIN
	result    <= sub_wire0(47 DOWNTO 0);

	lpm_xor_component : lpm_xor
	GENERIC MAP (
		lpm_size => 48,
		lpm_type => "LPM_XOR",
		lpm_width => 48
	)
	PORT MAP (
		data => data,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: CompactSymbol NUMERIC "0"
-- Retrieval info: PRIVATE: GateFunction NUMERIC "2"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: PRIVATE: InputAsBus NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WidthInput NUMERIC "48"
-- Retrieval info: PRIVATE: nInput NUMERIC "48"
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "48"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_XOR"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "48"
-- Retrieval info: USED_PORT: data 48 0 48 0 INPUT NODEFVAL data[47..0][47..0]
-- Retrieval info: USED_PORT: result 0 0 48 0 OUTPUT NODEFVAL result[47..0]
-- Retrieval info: CONNECT: @data 48 0 48 0 data 48 0 48 0
-- Retrieval info: CONNECT: result 0 0 48 0 @result 0 0 48 0
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL xor48.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL xor48.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL xor48.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL xor48.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL xor48_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
