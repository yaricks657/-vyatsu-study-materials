// megafunction wizard: %ALTFP_INV%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTFP_INV 

// ============================================================
// File Name: invert.v
// Megafunction Name(s):
// 			ALTFP_INV
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.1 Build 350 03/24/2010 SP 2 SJ Web Edition
// ************************************************************

//Copyright (C) 1991-2010 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module invert (
	clk_en,
	clock,
	data,
	result)/* synthesis synthesis_clearbox = 1 */;

	input	  clk_en;
	input	  clock;
	input	[46:0]  data;
	output	[46:0]  result;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_inv"
// Retrieval info: CONSTANT: PIPELINE NUMERIC "20"
// Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
// Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "11"
// Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "35"
// Retrieval info: USED_PORT: clk_en 0 0 0 0 INPUT NODEFVAL "clk_en"
// Retrieval info: CONNECT: @clk_en 0 0 0 0 clk_en 0 0 0 0
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: USED_PORT: data 0 0 47 0 INPUT NODEFVAL "data[46..0]"
// Retrieval info: CONNECT: @data 0 0 47 0 data 0 0 47 0
// Retrieval info: USED_PORT: result 0 0 47 0 OUTPUT NODEFVAL "result[46..0]"
// Retrieval info: CONNECT: result 0 0 47 0 @result 0 0 47 0
// Retrieval info: GEN_FILE: TYPE_NORMAL invert.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL invert.qip TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL invert.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL invert_inst.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL invert_bb.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL invert.inc TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL invert.cmp FALSE TRUE
// Retrieval info: LIB_FILE: lpm
